a::b.c
a #()::b.c
a::b#()::c.d
a # ( foo ) :: b # ( 1 ) :: c . d . e
