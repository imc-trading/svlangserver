[3:0]
abcd[1:0][2:0]
foo
bar [ 1:0 ]
