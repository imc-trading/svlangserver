"abcd"
""
"\\"
"\\\\"
"\\\\\\"
"\""
"\\\""
"\\\\\""
"\
\
"
